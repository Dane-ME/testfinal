module RISCV_Single_Cycle(
    input clk,
    input rst_n,
    output reg [31:0] PC,
    output wire [31:0] Inst
);
    wire [31:0] PC_next;
    wire [4:0] rs1, rs2, rd;
    wire [2:0] funct3;
    wire [6:0] opcode, funct7;
    wire [31:0] Imm;

    wire [31:0] ReadData1, ReadData2, WriteData;

    wire [31:0] ALU_in2, ALU_result;
    wire ALUZero;

    wire [31:0] MemReadData;

    wire [1:0] ALUSrc;
    wire [3:0] ALUCtrl;
    wire Branch, MemRead, MemWrite, MemToReg;
    wire RegWrite, PCSel;

    // PC update
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            PC <= 32'b0;
        else
            PC <= PC_next;
    end

    // Instruction Memory (IMEM)
    IMEM IMEM_inst(
        .addr(PC),
        .Instruction(Inst)
    );

    // Instruction field decoding
    assign opcode = Inst[6:0];
    assign rd     = Inst[11:7];
    assign funct3 = Inst[14:12];
    assign rs1    = Inst[19:15];
    assign rs2    = Inst[24:20];
    assign funct7 = Inst[31:25];

    // Immediate generator
    Imm_Gen imm_gen(
        .inst(Inst),
        .imm_out(Imm)
    );

    // Register File (instance name must be Reg_inst for tb)
    RegisterFile Reg_inst(
        .clk(clk),
        .rst_n(rst_n),
        .RegWrite(RegWrite),
        .rs1(rs1),
        .rs2(rs2),
        .rd(rd),
        .WriteData(WriteData),
        .ReadData1(ReadData1),
        .ReadData2(ReadData2)
    );

    // ALU input selection
    assign ALU_in2 = (ALUSrc[0]) ? Imm : ReadData2;

    // ALU
    ALU alu(
        .A(ReadData1),
        .B(ALU_in2),
        .ALUOp(ALUCtrl),
        .Result(ALU_result),
        .Zero(ALUZero)
    );

    // Data Memory (DMEM)
    DMEM DMEM_inst(
        .clk(clk),
        .rst_n(rst_n),
        .MemRead(MemRead),
        .MemWrite(MemWrite),
        .addr(ALU_result),
        .WriteData(ReadData2),
        .ReadData(MemReadData)
    );

    // Write-back mux
    assign WriteData = (MemToReg) ? MemReadData : ALU_result;

    // Control unit
    control_unit ctrl(
        .opcode(opcode),
        .funct3(funct3),
        .funct7(funct7),
        .ALUSrc(ALUSrc),
        .ALUOp(ALUCtrl),
        .Branch(Branch),
        .MemRead(MemRead),
        .MemWrite(MemWrite),
        .MemToReg(MemToReg),
        .RegWrite(RegWrite)
    );

    // Branch comparator
    Branch_Comp comp(
        .A(ReadData1),
        .B(ReadData2),
        .Branch(Branch),
        .funct3(funct3),
        .BrTaken(PCSel)
    );

    // Next PC logic
    assign PC_next = (PCSel) ? PC + Imm : PC + 4;

endmodule